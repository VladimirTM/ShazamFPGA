module twrom
(
input wire clk,
input wire twact,
input wire [10-1-2:0] twa,
output reg [16-1:0] twdr_cos
);


always @ ( posedge clk ) begin
if ( twact ) begin
case ( twa )
0: twdr_cos <= 32767;
1: twdr_cos <= 32766;
2: twdr_cos <= 32764;
3: twdr_cos <= 32761;
4: twdr_cos <= 32757;
5: twdr_cos <= 32751;
6: twdr_cos <= 32744;
7: twdr_cos <= 32736;
8: twdr_cos <= 32727;
9: twdr_cos <= 32717;
10: twdr_cos <= 32705;
11: twdr_cos <= 32692;
12: twdr_cos <= 32678;
13: twdr_cos <= 32662;
14: twdr_cos <= 32646;
15: twdr_cos <= 32628;
16: twdr_cos <= 32609;
17: twdr_cos <= 32588;
18: twdr_cos <= 32567;
19: twdr_cos <= 32544;
20: twdr_cos <= 32520;
21: twdr_cos <= 32495;
22: twdr_cos <= 32468;
23: twdr_cos <= 32441;
24: twdr_cos <= 32412;
25: twdr_cos <= 32382;
26: twdr_cos <= 32350;
27: twdr_cos <= 32318;
28: twdr_cos <= 32284;
29: twdr_cos <= 32249;
30: twdr_cos <= 32213;
31: twdr_cos <= 32175;
32: twdr_cos <= 32137;
33: twdr_cos <= 32097;
34: twdr_cos <= 32056;
35: twdr_cos <= 32014;
36: twdr_cos <= 31970;
37: twdr_cos <= 31926;
38: twdr_cos <= 31880;
39: twdr_cos <= 31833;
40: twdr_cos <= 31784;
41: twdr_cos <= 31735;
42: twdr_cos <= 31684;
43: twdr_cos <= 31633;
44: twdr_cos <= 31580;
45: twdr_cos <= 31525;
46: twdr_cos <= 31470;
47: twdr_cos <= 31413;
48: twdr_cos <= 31356;
49: twdr_cos <= 31297;
50: twdr_cos <= 31236;
51: twdr_cos <= 31175;
52: twdr_cos <= 31113;
53: twdr_cos <= 31049;
54: twdr_cos <= 30984;
55: twdr_cos <= 30918;
56: twdr_cos <= 30851;
57: twdr_cos <= 30783;
58: twdr_cos <= 30713;
59: twdr_cos <= 30643;
60: twdr_cos <= 30571;
61: twdr_cos <= 30498;
62: twdr_cos <= 30424;
63: twdr_cos <= 30349;
64: twdr_cos <= 30272;
65: twdr_cos <= 30195;
66: twdr_cos <= 30116;
67: twdr_cos <= 30036;
68: twdr_cos <= 29955;
69: twdr_cos <= 29873;
70: twdr_cos <= 29790;
71: twdr_cos <= 29706;
72: twdr_cos <= 29620;
73: twdr_cos <= 29534;
74: twdr_cos <= 29446;
75: twdr_cos <= 29358;
76: twdr_cos <= 29268;
77: twdr_cos <= 29177;
78: twdr_cos <= 29085;
79: twdr_cos <= 28992;
80: twdr_cos <= 28897;
81: twdr_cos <= 28802;
82: twdr_cos <= 28706;
83: twdr_cos <= 28608;
84: twdr_cos <= 28510;
85: twdr_cos <= 28410;
86: twdr_cos <= 28309;
87: twdr_cos <= 28207;
88: twdr_cos <= 28105;
89: twdr_cos <= 28001;
90: twdr_cos <= 27896;
91: twdr_cos <= 27790;
92: twdr_cos <= 27683;
93: twdr_cos <= 27575;
94: twdr_cos <= 27465;
95: twdr_cos <= 27355;
96: twdr_cos <= 27244;
97: twdr_cos <= 27132;
98: twdr_cos <= 27019;
99: twdr_cos <= 26904;
100: twdr_cos <= 26789;
101: twdr_cos <= 26673;
102: twdr_cos <= 26556;
103: twdr_cos <= 26437;
104: twdr_cos <= 26318;
105: twdr_cos <= 26198;
106: twdr_cos <= 26076;
107: twdr_cos <= 25954;
108: twdr_cos <= 25831;
109: twdr_cos <= 25707;
110: twdr_cos <= 25582;
111: twdr_cos <= 25456;
112: twdr_cos <= 25329;
113: twdr_cos <= 25200;
114: twdr_cos <= 25072;
115: twdr_cos <= 24942;
116: twdr_cos <= 24811;
117: twdr_cos <= 24679;
118: twdr_cos <= 24546;
119: twdr_cos <= 24413;
120: twdr_cos <= 24278;
121: twdr_cos <= 24143;
122: twdr_cos <= 24006;
123: twdr_cos <= 23869;
124: twdr_cos <= 23731;
125: twdr_cos <= 23592;
126: twdr_cos <= 23452;
127: twdr_cos <= 23311;
128: twdr_cos <= 23169;
129: twdr_cos <= 23026;
130: twdr_cos <= 22883;
131: twdr_cos <= 22739;
132: twdr_cos <= 22593;
133: twdr_cos <= 22447;
134: twdr_cos <= 22300;
135: twdr_cos <= 22153;
136: twdr_cos <= 22004;
137: twdr_cos <= 21855;
138: twdr_cos <= 21705;
139: twdr_cos <= 21554;
140: twdr_cos <= 21402;
141: twdr_cos <= 21249;
142: twdr_cos <= 21096;
143: twdr_cos <= 20941;
144: twdr_cos <= 20786;
145: twdr_cos <= 20630;
146: twdr_cos <= 20474;
147: twdr_cos <= 20317;
148: twdr_cos <= 20158;
149: twdr_cos <= 20000;
150: twdr_cos <= 19840;
151: twdr_cos <= 19680;
152: twdr_cos <= 19518;
153: twdr_cos <= 19357;
154: twdr_cos <= 19194;
155: twdr_cos <= 19031;
156: twdr_cos <= 18867;
157: twdr_cos <= 18702;
158: twdr_cos <= 18536;
159: twdr_cos <= 18370;
160: twdr_cos <= 18203;
161: twdr_cos <= 18036;
162: twdr_cos <= 17868;
163: twdr_cos <= 17699;
164: twdr_cos <= 17529;
165: twdr_cos <= 17359;
166: twdr_cos <= 17188;
167: twdr_cos <= 17017;
168: twdr_cos <= 16845;
169: twdr_cos <= 16672;
170: twdr_cos <= 16498;
171: twdr_cos <= 16324;
172: twdr_cos <= 16150;
173: twdr_cos <= 15975;
174: twdr_cos <= 15799;
175: twdr_cos <= 15622;
176: twdr_cos <= 15445;
177: twdr_cos <= 15268;
178: twdr_cos <= 15089;
179: twdr_cos <= 14911;
180: twdr_cos <= 14731;
181: twdr_cos <= 14551;
182: twdr_cos <= 14371;
183: twdr_cos <= 14190;
184: twdr_cos <= 14009;
185: twdr_cos <= 13827;
186: twdr_cos <= 13644;
187: twdr_cos <= 13461;
188: twdr_cos <= 13277;
189: twdr_cos <= 13093;
190: twdr_cos <= 12909;
191: twdr_cos <= 12724;
192: twdr_cos <= 12538;
193: twdr_cos <= 12352;
194: twdr_cos <= 12166;
195: twdr_cos <= 11979;
196: twdr_cos <= 11792;
197: twdr_cos <= 11604;
198: twdr_cos <= 11415;
199: twdr_cos <= 11227;
200: twdr_cos <= 11038;
201: twdr_cos <= 10848;
202: twdr_cos <= 10658;
203: twdr_cos <= 10468;
204: twdr_cos <= 10277;
205: twdr_cos <= 10086;
206: twdr_cos <= 9895;
207: twdr_cos <= 9703;
208: twdr_cos <= 9511;
209: twdr_cos <= 9318;
210: twdr_cos <= 9125;
211: twdr_cos <= 8932;
212: twdr_cos <= 8738;
213: twdr_cos <= 8544;
214: twdr_cos <= 8350;
215: twdr_cos <= 8155;
216: twdr_cos <= 7960;
217: twdr_cos <= 7765;
218: twdr_cos <= 7570;
219: twdr_cos <= 7374;
220: twdr_cos <= 7178;
221: twdr_cos <= 6982;
222: twdr_cos <= 6785;
223: twdr_cos <= 6588;
224: twdr_cos <= 6391;
225: twdr_cos <= 6194;
226: twdr_cos <= 5996;
227: twdr_cos <= 5799;
228: twdr_cos <= 5601;
229: twdr_cos <= 5402;
230: twdr_cos <= 5204;
231: twdr_cos <= 5005;
232: twdr_cos <= 4807;
233: twdr_cos <= 4608;
234: twdr_cos <= 4408;
235: twdr_cos <= 4209;
236: twdr_cos <= 4010;
237: twdr_cos <= 3810;
238: twdr_cos <= 3610;
239: twdr_cos <= 3410;
240: twdr_cos <= 3210;
241: twdr_cos <= 3010;
242: twdr_cos <= 2810;
243: twdr_cos <= 2610;
244: twdr_cos <= 2409;
245: twdr_cos <= 2209;
246: twdr_cos <= 2008;
247: twdr_cos <= 1807;
248: twdr_cos <= 1606;
249: twdr_cos <= 1406;
250: twdr_cos <= 1205;
251: twdr_cos <= 1004;
252: twdr_cos <= 803;
253: twdr_cos <= 602;
254: twdr_cos <= 401;
255: twdr_cos <= 200;
endcase
end
end
endmodule


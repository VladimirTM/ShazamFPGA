module twrom
(
input wire clk,
input wire twact,
input wire [10-1-2:0] twa,
output reg [15-1:0] twdr_cos
);


always @ ( posedge clk ) begin
if ( twact ) begin
case ( twa )
0: twdr_cos <= 16384;
1: twdr_cos <= 16384;
2: twdr_cos <= 16383;
3: twdr_cos <= 16381;
4: twdr_cos <= 16379;
5: twdr_cos <= 16376;
6: twdr_cos <= 16373;
7: twdr_cos <= 16369;
8: twdr_cos <= 16364;
9: twdr_cos <= 16359;
10: twdr_cos <= 16353;
11: twdr_cos <= 16347;
12: twdr_cos <= 16340;
13: twdr_cos <= 16332;
14: twdr_cos <= 16324;
15: twdr_cos <= 16315;
16: twdr_cos <= 16305;
17: twdr_cos <= 16295;
18: twdr_cos <= 16284;
19: twdr_cos <= 16273;
20: twdr_cos <= 16261;
21: twdr_cos <= 16248;
22: twdr_cos <= 16235;
23: twdr_cos <= 16221;
24: twdr_cos <= 16207;
25: twdr_cos <= 16192;
26: twdr_cos <= 16176;
27: twdr_cos <= 16160;
28: twdr_cos <= 16143;
29: twdr_cos <= 16125;
30: twdr_cos <= 16107;
31: twdr_cos <= 16088;
32: twdr_cos <= 16069;
33: twdr_cos <= 16049;
34: twdr_cos <= 16029;
35: twdr_cos <= 16008;
36: twdr_cos <= 15986;
37: twdr_cos <= 15964;
38: twdr_cos <= 15941;
39: twdr_cos <= 15917;
40: twdr_cos <= 15893;
41: twdr_cos <= 15868;
42: twdr_cos <= 15843;
43: twdr_cos <= 15817;
44: twdr_cos <= 15791;
45: twdr_cos <= 15763;
46: twdr_cos <= 15736;
47: twdr_cos <= 15707;
48: twdr_cos <= 15679;
49: twdr_cos <= 15649;
50: twdr_cos <= 15619;
51: twdr_cos <= 15588;
52: twdr_cos <= 15557;
53: twdr_cos <= 15525;
54: twdr_cos <= 15493;
55: twdr_cos <= 15460;
56: twdr_cos <= 15426;
57: twdr_cos <= 15392;
58: twdr_cos <= 15357;
59: twdr_cos <= 15322;
60: twdr_cos <= 15286;
61: twdr_cos <= 15250;
62: twdr_cos <= 15213;
63: twdr_cos <= 15175;
64: twdr_cos <= 15137;
65: twdr_cos <= 15098;
66: twdr_cos <= 15059;
67: twdr_cos <= 15019;
68: twdr_cos <= 14978;
69: twdr_cos <= 14937;
70: twdr_cos <= 14896;
71: twdr_cos <= 14854;
72: twdr_cos <= 14811;
73: twdr_cos <= 14768;
74: twdr_cos <= 14724;
75: twdr_cos <= 14680;
76: twdr_cos <= 14635;
77: twdr_cos <= 14589;
78: twdr_cos <= 14543;
79: twdr_cos <= 14497;
80: twdr_cos <= 14449;
81: twdr_cos <= 14402;
82: twdr_cos <= 14354;
83: twdr_cos <= 14305;
84: twdr_cos <= 14256;
85: twdr_cos <= 14206;
86: twdr_cos <= 14155;
87: twdr_cos <= 14104;
88: twdr_cos <= 14053;
89: twdr_cos <= 14001;
90: twdr_cos <= 13949;
91: twdr_cos <= 13896;
92: twdr_cos <= 13842;
93: twdr_cos <= 13788;
94: twdr_cos <= 13733;
95: twdr_cos <= 13678;
96: twdr_cos <= 13623;
97: twdr_cos <= 13567;
98: twdr_cos <= 13510;
99: twdr_cos <= 13453;
100: twdr_cos <= 13395;
101: twdr_cos <= 13337;
102: twdr_cos <= 13279;
103: twdr_cos <= 13219;
104: twdr_cos <= 13160;
105: twdr_cos <= 13100;
106: twdr_cos <= 13039;
107: twdr_cos <= 12978;
108: twdr_cos <= 12916;
109: twdr_cos <= 12854;
110: twdr_cos <= 12792;
111: twdr_cos <= 12729;
112: twdr_cos <= 12665;
113: twdr_cos <= 12601;
114: twdr_cos <= 12537;
115: twdr_cos <= 12472;
116: twdr_cos <= 12406;
117: twdr_cos <= 12340;
118: twdr_cos <= 12274;
119: twdr_cos <= 12207;
120: twdr_cos <= 12140;
121: twdr_cos <= 12072;
122: twdr_cos <= 12004;
123: twdr_cos <= 11935;
124: twdr_cos <= 11866;
125: twdr_cos <= 11797;
126: twdr_cos <= 11727;
127: twdr_cos <= 11656;
128: twdr_cos <= 11585;
129: twdr_cos <= 11514;
130: twdr_cos <= 11442;
131: twdr_cos <= 11370;
132: twdr_cos <= 11297;
133: twdr_cos <= 11224;
134: twdr_cos <= 11151;
135: twdr_cos <= 11077;
136: twdr_cos <= 11003;
137: twdr_cos <= 10928;
138: twdr_cos <= 10853;
139: twdr_cos <= 10778;
140: twdr_cos <= 10702;
141: twdr_cos <= 10625;
142: twdr_cos <= 10549;
143: twdr_cos <= 10471;
144: twdr_cos <= 10394;
145: twdr_cos <= 10316;
146: twdr_cos <= 10238;
147: twdr_cos <= 10159;
148: twdr_cos <= 10080;
149: twdr_cos <= 10001;
150: twdr_cos <= 9921;
151: twdr_cos <= 9841;
152: twdr_cos <= 9760;
153: twdr_cos <= 9679;
154: twdr_cos <= 9598;
155: twdr_cos <= 9516;
156: twdr_cos <= 9434;
157: twdr_cos <= 9352;
158: twdr_cos <= 9269;
159: twdr_cos <= 9186;
160: twdr_cos <= 9102;
161: twdr_cos <= 9019;
162: twdr_cos <= 8935;
163: twdr_cos <= 8850;
164: twdr_cos <= 8765;
165: twdr_cos <= 8680;
166: twdr_cos <= 8595;
167: twdr_cos <= 8509;
168: twdr_cos <= 8423;
169: twdr_cos <= 8337;
170: twdr_cos <= 8250;
171: twdr_cos <= 8163;
172: twdr_cos <= 8076;
173: twdr_cos <= 7988;
174: twdr_cos <= 7900;
175: twdr_cos <= 7812;
176: twdr_cos <= 7723;
177: twdr_cos <= 7635;
178: twdr_cos <= 7545;
179: twdr_cos <= 7456;
180: twdr_cos <= 7366;
181: twdr_cos <= 7276;
182: twdr_cos <= 7186;
183: twdr_cos <= 7096;
184: twdr_cos <= 7005;
185: twdr_cos <= 6914;
186: twdr_cos <= 6823;
187: twdr_cos <= 6731;
188: twdr_cos <= 6639;
189: twdr_cos <= 6547;
190: twdr_cos <= 6455;
191: twdr_cos <= 6363;
192: twdr_cos <= 6270;
193: twdr_cos <= 6177;
194: twdr_cos <= 6084;
195: twdr_cos <= 5990;
196: twdr_cos <= 5897;
197: twdr_cos <= 5803;
198: twdr_cos <= 5708;
199: twdr_cos <= 5614;
200: twdr_cos <= 5520;
201: twdr_cos <= 5425;
202: twdr_cos <= 5330;
203: twdr_cos <= 5235;
204: twdr_cos <= 5139;
205: twdr_cos <= 5044;
206: twdr_cos <= 4948;
207: twdr_cos <= 4852;
208: twdr_cos <= 4756;
209: twdr_cos <= 4660;
210: twdr_cos <= 4563;
211: twdr_cos <= 4467;
212: twdr_cos <= 4370;
213: twdr_cos <= 4273;
214: twdr_cos <= 4176;
215: twdr_cos <= 4078;
216: twdr_cos <= 3981;
217: twdr_cos <= 3883;
218: twdr_cos <= 3786;
219: twdr_cos <= 3688;
220: twdr_cos <= 3590;
221: twdr_cos <= 3492;
222: twdr_cos <= 3393;
223: twdr_cos <= 3295;
224: twdr_cos <= 3196;
225: twdr_cos <= 3098;
226: twdr_cos <= 2999;
227: twdr_cos <= 2900;
228: twdr_cos <= 2801;
229: twdr_cos <= 2702;
230: twdr_cos <= 2603;
231: twdr_cos <= 2503;
232: twdr_cos <= 2404;
233: twdr_cos <= 2305;
234: twdr_cos <= 2205;
235: twdr_cos <= 2105;
236: twdr_cos <= 2006;
237: twdr_cos <= 1906;
238: twdr_cos <= 1806;
239: twdr_cos <= 1706;
240: twdr_cos <= 1606;
241: twdr_cos <= 1506;
242: twdr_cos <= 1406;
243: twdr_cos <= 1306;
244: twdr_cos <= 1205;
245: twdr_cos <= 1105;
246: twdr_cos <= 1005;
247: twdr_cos <= 904;
248: twdr_cos <= 804;
249: twdr_cos <= 704;
250: twdr_cos <= 603;
251: twdr_cos <= 503;
252: twdr_cos <= 402;
253: twdr_cos <= 302;
254: twdr_cos <= 201;
255: twdr_cos <= 101;
endcase
end
end
endmodule

